library verilog;
use verilog.vl_types.all;
entity TN4_vlg_vec_tst is
end TN4_vlg_vec_tst;
