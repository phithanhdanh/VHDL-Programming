library verilog;
use verilog.vl_types.all;
entity TN4_Behavioral_vlg_vec_tst is
end TN4_Behavioral_vlg_vec_tst;
