library verilog;
use verilog.vl_types.all;
entity TN5_vlg_vec_tst is
end TN5_vlg_vec_tst;
